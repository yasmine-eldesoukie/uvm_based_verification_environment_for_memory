package mem_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    `include "interface.sv"

    import seq_item_pkg::*;
    import driver_pkg::*;
	import monitor_pkg::*;
	import sequencer_pkg::*;
	import agent_pkg::*;
	import scoreboard_pkg::*;
	import subscriber_pkg::*;
	import env_pkg::*;
	import sequence_pkg::*;
	import test_pkg::*;
endpackage