package driver_pkg;
	class my_driver extends uvm_driver #(my_seq_item);

    endclass
endpackage

