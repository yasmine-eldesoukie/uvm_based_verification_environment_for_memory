package sequencer_pkg;
	class my_sequencer extends uvm_sequencer #(my_seq_item);

    endclass
endpackage
