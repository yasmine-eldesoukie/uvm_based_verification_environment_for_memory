package env_pkg;
	class my_env extends uvm_env;

    endclass
endpackage
