package seq_item_pkg;
    class my_seq_item extends uvm_sequence_item;
            
    endclass
endpackage
