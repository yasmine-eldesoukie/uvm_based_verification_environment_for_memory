package agent_pkg;
	class my_agent extends uvm_agent;

    endclass
endpackage
