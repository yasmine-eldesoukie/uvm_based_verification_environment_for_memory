package scoreborad_pkg;
	class my_scoreborad extends uvm_scoreborad #(my_seq_item);

    endclass
endpackage
