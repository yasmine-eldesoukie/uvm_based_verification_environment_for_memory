package test_pkg;
	class my_test extends uvm_test;

    endclass
endpackage
