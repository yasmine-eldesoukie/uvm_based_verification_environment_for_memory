package monitor_pkg;
	class my_monitor extends uvm_monitor;

    endclass
endpackage
