package sequence_pkg;
	class my_sequence extends uvm_sequence #(my_seq_item);

    endclass
endpackage
